`timescale 1ns / 1ps

module SPHY_Wave_Generator (
    input wire clk,           // High-speed system clock
    input wire reset,         // Active-high reset
    input wire [11:0] feedback_in, // From ADC (Infinite Loop Feedback)
    output reg [11:0] hphyspi,// Primary harmonic stabilizer wave amplitude
    output reg [11:0] sphyspi // Secondary phase-alignment wave amplitude
);
    // Phase accumulators to track the current position in the wave cycle
    reg [23:0] phase_acc_h;
    reg [23:0] phase_acc_s;
    
    // Tuning parameters for the wave frequencies
    parameter FREQ_H = 24'd419430; 
    parameter FREQ_S = 24'd838860; 
    
    // Look-Up Table (LUT) holding the pre-calculated SPHY wave geometry
    reg [11:0] sphy_lut [0:255];
    
    // Load the wave memory file generated by the Q-OS Python engine
    initial $readmemh("sphy_table.mem", sphy_lut);

    always @(posedge clk) begin
        if (reset) begin
            phase_acc_h <= 24'd0;
            phase_acc_s <= 24'd0;
            hphyspi <= 12'd0;
            sphyspi <= 12'd0;
        end else begin
            // INFINITE LOOP MODULATION:
            // The feedback_in (ADC value) modulates the phase accumulation speed.
            // This creates the 'Phase-Locked' behavior described in v2.0.
            // We shift feedback up to have a significant effect on the 24-bit accumulator.
            phase_acc_h <= phase_acc_h + FREQ_H + {feedback_in, 4'b0};
            phase_acc_s <= phase_acc_s + FREQ_S + {feedback_in, 4'b0};
            
            // Map the top 8 bits of the accumulator to the 256-value LUT
            hphyspi <= sphy_lut[phase_acc_h[23:16]];
            sphyspi <= sphy_lut[phase_acc_s[23:16]];
        end
    end
endmodule